`timescale 1ns / 1ps

module TopMicro(
    input [15:0] sw,
    input btnC,
    input clk,
    output [15:0] led
);

    reg clkdiv = 0;
    integer i = 0;

    localparam st_Idle = 0;
    localparam st_Presionado = 1;

    reg [1:0] estado = st_Idle;

    always @( posedge clk ) begin

        case (estado)

            st_Idle: begin
                if (btnC == 1) estado <= st_Presionado;
                clkdiv <= 0;
            end

            st_Presionado: begin
                clkdiv <= 1;
                if ( i < 50_000_000 ) i = i + 1;
                else begin
                    i = 0;
                    estado <= st_Idle;
                end
            end

        endcase
    end

    // 1111_1111_1111_0111_0000_0000_0000_0010
    // 1111_1111_1111_0111_0000_0000_0000_0001
    // 0000_0000_0000_1000_1111_1111_1111_1110
    
    // 3128_2724_2320_1916_1512_1108_0704_0300
    // 1000_0000_0010_0111_0000_0000_0110_1111
    // 1111_1111_1111_0111_0000_0000_0000_0010
    //                1000_1111_1111_1111_1110
    //                                   8FFFE



    // 1000_0000_0010_0111_0000_0000_0110_1111
    // 1111_1111_1011_1111_1111_0000_0110_1111
    // FFBFF06F
    // -6 = 1010 = 1111_1111_1111_1111_1101

    //
    //
    // -6 = 0110 -> 111111010, entonces necesitamos escribir un 1111_1111_1111_1111_1101 -> 1111100 -> 000011
    // FFFF_FFFD

    // 2017_1613_1209_0805_0401
    // 1111_1111_1111_1111_1101
    // 1.11_1111_1101.1.111_1111_1._0000_0110_1111
    // 1111_1111_1011_1111_1111_0000_0110_1111
    // FFBFF06F

    // -6*4 = -24 = -01_1000 =
    // 
    // 2017_1613_1209_0805_0401
    // 1111_1111_1111_1110_1000
    // 1.11_1110_1000.1.111_1111_1.00000.1101111
    // 1111_1101_0001_1111_1111_0000_0110_1111
    // FB1FF06F -> fb1ff06f

    // -6*4 = -24 = -01_1000 =
    // 
    // 2017_1613_1209_0805_0401
    // 1111_1111_1111_1111_0100
    // 1.11_1111_0100.1.111_1111_1.00000.1101111
    // 1111_1110_1001_1111_1111_0000_0110_1111
    // FE6FF06F -> fe6ff06f
        
    //       |func7 ||rs2 | |rs1 ||3| |rd  ||opcode|
    reg [32 * 12 - 1:0] instruction_bank = {           //
        {32'b1111_1111_1011_1111_1111_0000_0110_1111}, //  0000_0000_0000_0101_1000_0100_0110_0011 
        {32'b0000_0000_0001_0000_0000_0010_0001_0011}, //
        {32'b0000_0000_0001_0001_1111_0010_0001_0011}, // 
        {32'b0000_0000_0011_0000_0010_0000_1000_0011}, //
        {32'b0000_0000_1010_0000_1111_0001_0001_0011}, //
        {32'b0000_0000_0010_0000_0010_0001_1010_0011}, //
        {32'b1111_1110_0000_0000_1000_1110_1110_0011}, //
        {32'b1111_1111_0001_1111_1111_0000_0110_1111}, //
        {32'b1010_1001_1010_1011_1010_1010_1010_1010}, //
        {32'b1010_1001_1010_1011_1010_1010_1010_1010}, //
        {32'b1010_1001_1010_1011_1010_1010_1010_1010}, //
        {32'b1010_1001_1010_1011_1010_1010_1010_1010}  //
    };

    wire reset;
    wire [31:0] Progin;
    wire [31:0] Datain;
    wire [31:0] Progaddress;
    wire WE;
    wire [31:0] address;
    wire [31:0] Dataout;
    wire [31:0] i_debug;
    wire [31:0] o_debug;

    assign reset = sw[15];
    assign Progin = instruction_bank[((12-1)*4-Progaddress)*8 +: 32];
    // assign Datain = 32'b0 | sw[3:0];

    assign i_debug[15:0] = sw[15:0];
    assign led[15:0] = address[15:0];//o_debug[15:0];
    // assign led[2:0] = o_debug[2:0];
    // assign led[5:3] = Dataout[3:0];
    // assign led[9:6] = address[3:0];
    // assign led[14:10] = Progaddress[4:0];
    // assign led[15] = WE;

    Microprocesador micro (
        clkdiv,
        reset,
        Progin,
        Datain,
        Progaddress,
        WE,
        address,
        Dataout,
        i_debug,
        o_debug
    );

    // assign led = debug[15:0];

endmodule