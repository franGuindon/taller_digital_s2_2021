`timescale 1ns / 1ps

module CLA_4bit(output [3:0] S,
		output 	     Cout,
		input [3:0]  A,B,
		input 	     Cin);
   
   wire [3:0] 		     G,P,C;
   
   assign G = A & B; //Generate
   assign P = A ^ B; //Propagate
   assign C[0] = Cin;
   assign C[1] = G[0] | (P[0] & C[0]);
   assign C[2] = G[1] | (P[1] & G[0]) | (P[1] & P[0] & C[0]);
   assign C[3] = G[2] | (P[2] & G[1]) | (P[2] & P[1] & G[0]) | (P[2] & P[1] & P[0] & C[0]);
   assign Cout = G[3] | (P[3] & G[2]) | (P[3] & P[2] & G[1]) | (P[3] & P[2] & P[1] & G[0]) |(P[3] & P[2] & P[1] & P[0] & C[0]);
   assign S = P ^ C;
   
endmodule
